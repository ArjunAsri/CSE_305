LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_SIGNED.all;

ENTITY ONE_SECOND_CLOCK IS 
PORT ( SIGNAl CLOCK 			:IN STD_LOGIC;
		 SIGNAL CLOCK_OUT : OUT STD_LOGIC;
		 SIGNAL ENABLE_OUT : OUT STD_LOGIC );
END ONE_SECOND_CLOCK;


ARCHITECTURE BEHAVIOUR OF ONE_SECOND_CLOCK IS

-- SIGNAL t_BULLET_X_POSITION : STD_LOGIC_VECTOR (10 DOWNTO 0) := '0' & MOUSE_COLUMN;
SIGNAL CLOCK_STATE : STD_LOGIC := '0';
BEGIN
 
PROCESS(CLOCK)
VARIABLE COUNTER : INTEGER RANGE 0 TO 12499999 := 0;
BEGIN

IF(RISING_EDGE(CLOCK)) THEN
	IF(COUNTER = 12499999)THEN
	COUNTER := 0;
	CLOCK_STATE <= '1';
	ELSE
	CLOCK_STATE <= '0';
	COUNTER := COUNTER +1;
	END IF;
-- THIS resets the enable to 0 and so now the player waits for fire signal
END IF;
END PROCESS;
CLOCK_OUT <= CLOCK_STATE;
END BEHAVIOUR;